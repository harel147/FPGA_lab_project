//-- Alex Grinshpun Apr 2017
//-- Dudy Nov 13 2017
// System-Verilog Alex Grinshpun May 2018
// New coding convention dudy December 2018
// (c) Technion IIT, Department of Electrical Engineering  May 2019 

module	objects_mux_all	(
//		--------	Clock Input		
					input		logic	clk,
					input		logic	resetN,
		// smiley 
					input		logic	smileyDrawingRequest, // two set of inputs per unit
					input		logic	[7:0] smileyRGB, 
		//square
					input		logic	squareDrawingRequest, // two set of inputs per unit
					input		logic	[7:0] squareRGB, 
		
		// background 
					input		logic	[7:0] backGroundRGB, 
		// add the box here 
					
				// fill your code here - inputs for box
					
					output	logic	[7:0] redOut, // full 24 bits color output
					output	logic	[7:0] greenOut, 
					output	logic	[7:0] blueOut 
);

logic [7:0] tmpRGB;


assign redOut	  = {tmpRGB[7:5], {5{tmpRGB[5]}}}; //--  extend LSB to create 10 bits per color  
assign greenOut  = {tmpRGB[4:2], {5{tmpRGB[2]}}};
assign blueOut	  = {tmpRGB[1:0], {6{tmpRGB[0]}}};

//======--------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
			tmpRGB	<= 8'b0;
	end
	else begin
		if (smileyDrawingRequest == 1'b1 )   
			tmpRGB <= smileyRGB;  //first priority 
		
		// fill your code here logics for box
		
		else if (squareDrawingRequest == 1'b1 )   
			tmpRGB <= squareRGB;  //second priority 
		
		// fill your code here logics for box
		
			else
			tmpRGB <= backGroundRGB ; // last priority 
		end ; 
	end

endmodule


